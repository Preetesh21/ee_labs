*Transmission Line 10 section with open ckt
V1 1 0 sin(0 20v 1.5khz)
R1 1 2 5
L1 2 3 2m
C1 3 0 0.47u
R2 3 0 1e4
R3 3 4 5
L2 4 5 2m
R4 5 6 5
L3 6 7  2m
C2 7 0 0.47u
R5 7 0 1e4
R6 7 8 5
L4 8 9 2m
R7 9 10 5
L5 10 11 2m
C3 11 0 0.47u
R8 11 0 1e4
R9 11 12 5
L6 12 13 2m
R10 13 14 5
L7 14 15 2m
C4 15 0 0.47u
R11 15 0 1e4
R12 15 16 5
L8 16 17 2m
R13 17 18 5
L9 18 19 2m
C5 19 0 0.47u
R14 19 0 1e4
R15 19 20 5
L10 20 21 2m
R16 21 22 5
L11 22 23 2m
C6 23 0 0.47u
R17 23 0 1e4
R18 23 24 5
L12 24 25 2m
R19 25 26 5
L13 26 27 2m
C7 27 0 0.47u
R20 27 0 1e4
R21 27 28 5
L14 28 29 2m
R22 29 30 5
L15 30 31 2m
C8 31 0 0.47u
R23 31 0 1e4
R24 31 32 5
L16 32 33 2m
R25 33 34 5
L17 34 35 2m
C9 35 0 0.47u
R26 35 0 1e4
R27 35 36 5
L18 36 37 2m
R28 37 38 5
L19 38 39 2m
C10 39 0 0.47u
R29 39 0 1e4
R30 39 40 5
L20 40 41 2m
R36 41 0 93.37
.tran 0 10ms [0 100ns]
.probe